`timescale 10ns/1ps
module andgate(a,b,y);
input a,b;
output y;

assign z= a&b;

endmodule
